//                              -*- Mode: Verilog -*-
// Filename        : foo.v
// Description     : GIT TESTING
// Author          : Phil Tracton
// Created On      : Mon Feb 20 21:46:47 2012
// Last Modified By: .
// Last Modified On: .
// Update Count    : 0
// Status          : Unknown, Use with caution!


module foo(input wire clk,
	   input wire rst,
	   input wire rx,
	   output reg tx
	   );


endmodule // foo
